`define CONNECT signals_if(.data_out[0][0][0](DUT._rw_[1]._clm_[1].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[0][0][0](DUT._rw_[1]._clm_[1].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][0][1](DUT._rw_[1]._clm_[1].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[0][0][1](DUT._rw_[1]._clm_[1].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][0][2](DUT._rw_[1]._clm_[1].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[0][0][2](DUT._rw_[1]._clm_[1].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][0][3](DUT._rw_[1]._clm_[1].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[0][0][3](DUT._rw_[1]._clm_[1].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][1][0](DUT._rw_[1]._clm_[2].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[0][1][0](DUT._rw_[1]._clm_[2].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][1][1](DUT._rw_[1]._clm_[2].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[0][1][1](DUT._rw_[1]._clm_[2].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][1][2](DUT._rw_[1]._clm_[2].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[0][1][2](DUT._rw_[1]._clm_[2].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][1][3](DUT._rw_[1]._clm_[2].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[0][1][3](DUT._rw_[1]._clm_[2].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][2][0](DUT._rw_[1]._clm_[3].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[0][2][0](DUT._rw_[1]._clm_[3].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][2][1](DUT._rw_[1]._clm_[3].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[0][2][1](DUT._rw_[1]._clm_[3].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][2][2](DUT._rw_[1]._clm_[3].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[0][2][2](DUT._rw_[1]._clm_[3].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][2][3](DUT._rw_[1]._clm_[3].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[0][2][3](DUT._rw_[1]._clm_[3].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][3][0](DUT._rw_[1]._clm_[4].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[0][3][0](DUT._rw_[1]._clm_[4].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][3][1](DUT._rw_[1]._clm_[4].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[0][3][1](DUT._rw_[1]._clm_[4].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][3][2](DUT._rw_[1]._clm_[4].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[0][3][2](DUT._rw_[1]._clm_[4].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[0][3][3](DUT._rw_[1]._clm_[4].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[0][3][3](DUT._rw_[1]._clm_[4].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][0][0](DUT._rw_[2]._clm_[1].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[1][0][0](DUT._rw_[2]._clm_[1].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][0][1](DUT._rw_[2]._clm_[1].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[1][0][1](DUT._rw_[2]._clm_[1].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][0][2](DUT._rw_[2]._clm_[1].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[1][0][2](DUT._rw_[2]._clm_[1].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][0][3](DUT._rw_[2]._clm_[1].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[1][0][3](DUT._rw_[2]._clm_[1].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][1][0](DUT._rw_[2]._clm_[2].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[1][1][0](DUT._rw_[2]._clm_[2].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][1][1](DUT._rw_[2]._clm_[2].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[1][1][1](DUT._rw_[2]._clm_[2].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][1][2](DUT._rw_[2]._clm_[2].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[1][1][2](DUT._rw_[2]._clm_[2].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][1][3](DUT._rw_[2]._clm_[2].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[1][1][3](DUT._rw_[2]._clm_[2].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][2][0](DUT._rw_[2]._clm_[3].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[1][2][0](DUT._rw_[2]._clm_[3].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][2][1](DUT._rw_[2]._clm_[3].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[1][2][1](DUT._rw_[2]._clm_[3].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][2][2](DUT._rw_[2]._clm_[3].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[1][2][2](DUT._rw_[2]._clm_[3].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][2][3](DUT._rw_[2]._clm_[3].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[1][2][3](DUT._rw_[2]._clm_[3].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][3][0](DUT._rw_[2]._clm_[4].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[1][3][0](DUT._rw_[2]._clm_[4].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][3][1](DUT._rw_[2]._clm_[4].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[1][3][1](DUT._rw_[2]._clm_[4].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][3][2](DUT._rw_[2]._clm_[4].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[1][3][2](DUT._rw_[2]._clm_[4].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[1][3][3](DUT._rw_[2]._clm_[4].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[1][3][3](DUT._rw_[2]._clm_[4].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][0][0](DUT._rw_[3]._clm_[1].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[2][0][0](DUT._rw_[3]._clm_[1].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][0][1](DUT._rw_[3]._clm_[1].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[2][0][1](DUT._rw_[3]._clm_[1].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][0][2](DUT._rw_[3]._clm_[1].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[2][0][2](DUT._rw_[3]._clm_[1].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][0][3](DUT._rw_[3]._clm_[1].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[2][0][3](DUT._rw_[3]._clm_[1].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][1][0](DUT._rw_[3]._clm_[2].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[2][1][0](DUT._rw_[3]._clm_[2].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][1][1](DUT._rw_[3]._clm_[2].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[2][1][1](DUT._rw_[3]._clm_[2].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][1][2](DUT._rw_[3]._clm_[2].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[2][1][2](DUT._rw_[3]._clm_[2].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][1][3](DUT._rw_[3]._clm_[2].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[2][1][3](DUT._rw_[3]._clm_[2].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][2][0](DUT._rw_[3]._clm_[3].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[2][2][0](DUT._rw_[3]._clm_[3].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][2][1](DUT._rw_[3]._clm_[3].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[2][2][1](DUT._rw_[3]._clm_[3].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][2][2](DUT._rw_[3]._clm_[3].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[2][2][2](DUT._rw_[3]._clm_[3].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][2][3](DUT._rw_[3]._clm_[3].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[2][2][3](DUT._rw_[3]._clm_[3].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][3][0](DUT._rw_[3]._clm_[4].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[2][3][0](DUT._rw_[3]._clm_[4].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][3][1](DUT._rw_[3]._clm_[4].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[2][3][1](DUT._rw_[3]._clm_[4].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][3][2](DUT._rw_[3]._clm_[4].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[2][3][2](DUT._rw_[3]._clm_[4].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[2][3][3](DUT._rw_[3]._clm_[4].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[2][3][3](DUT._rw_[3]._clm_[4].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][0][0](DUT._rw_[4]._clm_[1].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[3][0][0](DUT._rw_[4]._clm_[1].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][0][1](DUT._rw_[4]._clm_[1].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[3][0][1](DUT._rw_[4]._clm_[1].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][0][2](DUT._rw_[4]._clm_[1].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[3][0][2](DUT._rw_[4]._clm_[1].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][0][3](DUT._rw_[4]._clm_[1].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[3][0][3](DUT._rw_[4]._clm_[1].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][1][0](DUT._rw_[4]._clm_[2].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[3][1][0](DUT._rw_[4]._clm_[2].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][1][1](DUT._rw_[4]._clm_[2].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[3][1][1](DUT._rw_[4]._clm_[2].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][1][2](DUT._rw_[4]._clm_[2].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[3][1][2](DUT._rw_[4]._clm_[2].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][1][3](DUT._rw_[4]._clm_[2].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[3][1][3](DUT._rw_[4]._clm_[2].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][2][0](DUT._rw_[4]._clm_[3].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[3][2][0](DUT._rw_[4]._clm_[3].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][2][1](DUT._rw_[4]._clm_[3].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[3][2][1](DUT._rw_[4]._clm_[3].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][2][2](DUT._rw_[4]._clm_[3].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[3][2][2](DUT._rw_[4]._clm_[3].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][2][3](DUT._rw_[4]._clm_[3].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[3][2][3](DUT._rw_[4]._clm_[3].rtr._nu_[3].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][3][0](DUT._rw_[4]._clm_[4].rtr._nu_[0].rtr_ntrfs_.data_out), .pop[3][3][0](DUT._rw_[4]._clm_[4].rtr._nu_[0].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][3][1](DUT._rw_[4]._clm_[4].rtr._nu_[1].rtr_ntrfs_.data_out), .pop[3][3][1](DUT._rw_[4]._clm_[4].rtr._nu_[1].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][3][2](DUT._rw_[4]._clm_[4].rtr._nu_[2].rtr_ntrfs_.data_out), .pop[3][3][2](DUT._rw_[4]._clm_[4].rtr._nu_[2].rtr_ntrfs_.pop));  \
signals_if(.data_out[3][3][3](DUT._rw_[4]._clm_[4].rtr._nu_[3].rtr_ntrfs_.data_out), .pop[3][3][3](DUT._rw_[4]._clm_[4].rtr._nu_[3].rtr_ntrfs_.pop));
