class checker_scoreboard;
  ag_chk_sb_mbx ag_chk_sb_mbx;
  ag_chk_sb	ag_chk_sb_transaction;
  
  
  function new();
    
  endfunction 
  
  
  
endclass